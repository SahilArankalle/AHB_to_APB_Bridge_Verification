module top;

    import test_pkg::*;
    import uvm_pkg::*;


    initial
        begin
            run_test();
    
        end

endmodule
